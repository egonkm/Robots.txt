User-agent: *
Disallow: /HOME/
Disallow: /proxyDevice
Disallow: /proxydevice
Disallow: /gz/webdevice/config

