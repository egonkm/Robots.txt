#Build version: R718d
#Generated on: Fri May 24 01:00:00 EDT 2024

User-agent: *
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /flights/$
Allow: /hotels/$
Allow: /cars/$
Allow: /trains/$
Allow: /trips/users/
Allow: /cruises/$
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /charm/g/
Allow: /tweb/app/
Allow: /s/horizon/compareTo
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /api/search/V8
Allow: /charm/
Allow: /trips/$
Allow: /things-to-do/$
Disallow: /things-to-do/*
Disallow: /charm/horizon/cars/citycars/CityCarsAgencyMapViewLink
Disallow: /charm/horizon/cars/airportcars/AirportCarsResults
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /s/horizon/common/layout/StyleJamNavMenu
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/flights/flightdeals/frontdoor/FlightDealsLinks
Disallow: /charm/horizon/common/compareto/slide/SlideCompareToAction
Disallow: /charm/horizon/common/layout/MoreNavContentApiAction
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/flightroutes/AjaxGoodToKnow
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/flights/flightroutes/AjaxWhenToBookCharts
Disallow: /charm/horizon/flights/flightroutes/AjaxFlightRouteInfoTable
Disallow: /charm/horizon/flights/flightroutes/CountryCityRouteFAQAction
Disallow: /charm/horizon/flights/flightroutes/TravelRestrictionsNeededDocumentsFaqAction
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/common/upgrade/UpgradeBrowser
Disallow: /charm/horizon/flights/airport/AirportFlightStatusTable
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /s/horizon/common/corporate/PlatformToBusiness
Disallow: /charm/horizon/cars/citycars/CityCarsAgencyMap
Disallow: /charm/horizon/flights/airport/AirportMap
Disallow: /charm/horizon/flights/search/NonstopAvailabilityAction
Disallow: /vs/
Disallow: /%20/
Disallow: /maps/
Disallow: /tweb/
Disallow: /sem/
Disallow: /horizon/sem/
Disallow: /*/landing/*.html
Disallow: /semi/
Disallow: /hotels/
Disallow: /flights/
Disallow: /cars/
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /splitbookingflightreservation
Disallow: /splitbookinghotelreservation
Disallow: /book
Disallow: /rentals/
Disallow: /global
Disallow: /trains/
Disallow: /cruises/
Disallow: /huddle/
Disallow: /guides/u/*
Disallow: /guides/admin*
Disallow: /guides/missing
Disallow: /guides/noaccess
Disallow: /s/horizon/common/personalization/guidebooks/
Disallow: /restaurants/
Disallow: /ugtm
Disallow: /curated/
Disallow: /nearby/
Disallow: /platform2business
Disallow: /playground
Disallow: /sandbox
Disallow: /benchmark
Disallow: /charm/horizon/common/layout/SocialMediaLinks
Disallow: /charm/horizon/
Disallow: /nox/
Disallow: /gtm
Disallow: /mgtm
Disallow: /trips/
Disallow: /book/
Disallow: /picasso/place
Disallow: /charm/horizon/flights/flightroutes/AjaxPackageSearchForm
Disallow: /charm/horizon/hotels/cityguides/AjaxSeoCityGuidesFlightSearchForm
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/dynamicfrontdoor/v1/
Disallow: /mvm
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic
Disallow: /cimg/
Disallow: /in
Disallow: /news/search/

User-agent: Facebot
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /flights/$
Allow: /hotels/$
Allow: /cars/$
Allow: /trains/$
Allow: /trips/users/
Allow: /cruises/$
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /book
Allow: /charm/g/
Allow: /tweb/app/
Allow: /s/horizon/compareTo
Disallow: /charm/horizon/cars/citycars/CityCarsAgencyMapViewLink
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /s/horizon/common/layout/StyleJamNavMenu
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/flightroutes/AjaxGoodToKnow
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/flights/flightroutes/AjaxWhenToBookCharts
Disallow: /charm/horizon/flights/flightroutes/AjaxFlightRouteInfoTable
Disallow: /charm/horizon/flights/flightroutes/CountryCityRouteFAQAction
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /vs/
Disallow: /%20/
Disallow: /maps/
Disallow: /tweb/
Disallow: /sem/
Disallow: /horizon/sem/
Disallow: /*/landing/*.html
Disallow: /semi/
Disallow: /hotels/
Disallow: /flights/
Disallow: /cars/
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /splitbookingflightreservation
Disallow: /splitbookinghotelreservation
Disallow: /in
Disallow: /rentals/
Disallow: /trains/
Disallow: /cruises/
Disallow: /huddle/
Disallow: /guides/u/*
Disallow: /guides/admin*
Disallow: /guides/missing
Disallow: /guides/noaccess
Disallow: /s/horizon/common/personalization/guidebooks/
Disallow: /curated/
Disallow: /charm/horizon/flights/flightroutes/AjaxPackageSearchForm
Disallow: /charm/horizon/hotels/cityguides/AjaxSeoCityGuidesFlightSearchForm
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/dynamicfrontdoor/v1/
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic

User-agent: Twitterbot
Allow: /guides/u/*
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /flights/$
Allow: /hotels/$
Allow: /cars/$
Allow: /trains/$
Allow: /trips/users/
Allow: /cruises/$
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /book
Allow: /charm/g/
Allow: /tweb/app/
Allow: /s/horizon/compareTo
Disallow: /charm/horizon/cars/citycars/CityCarsAgencyMapViewLink
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /s/horizon/common/layout/StyleJamNavMenu
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/flightroutes/AjaxGoodToKnow
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/flights/flightroutes/AjaxWhenToBookCharts
Disallow: /charm/horizon/flights/flightroutes/AjaxFlightRouteInfoTable
Disallow: /charm/horizon/flights/flightroutes/CountryCityRouteFAQAction
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /vs/
Disallow: /%20/
Disallow: /maps/
Disallow: /tweb/
Disallow: /sem/
Disallow: /horizon/sem/
Disallow: /*/landing/*.html
Disallow: /semi/
Disallow: /hotels/
Disallow: /flights/
Disallow: /cars/
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /splitbookingflightreservation
Disallow: /splitbookinghotelreservation
Disallow: /in
Disallow: /rentals/
Disallow: /trains/
Disallow: /cruises/
Disallow: /huddle/
Disallow: /guides/admin*
Disallow: /guides/missing
Disallow: /guides/noaccess
Disallow: /s/horizon/common/personalization/guidebooks/
Disallow: /curated/
Disallow: /charm/horizon/flights/flightroutes/AjaxPackageSearchForm
Disallow: /charm/horizon/hotels/cityguides/AjaxSeoCityGuidesFlightSearchForm
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/dynamicfrontdoor/v1/
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic

User-agent: ChatGPT-User
Allow: /flights/
Allow: /hotels/
Allow: /cars/
Allow: /explore/
Allow: /sherlock/
Disallow: /api/
Disallow: /a/
Disallow: /i/
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /in
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/

User-agent: AdsBot-Google
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /api/search/V8
Allow: /tweb/hotels/results-ajax
Allow: /tweb/hotel/history/
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /hotels/$
Allow: /hotels/*
Allow: /flights/$
Allow: /flights/*
Allow: /cars/$
Allow: /cars/*
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /sem/
Allow: /semi/
Allow: /in
Allow: /horizon/sem/
Allow: /*/landing/*.html
Allow: /tweb/hotels/
Allow: /tweb/flights/
Allow: /tweb/cars/
Allow: /charm/
Allow: /book
Allow: /s/horizon/compareTo
Allow: /s/tweb/session/refresh/presentation
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/flights/airport/AirportFlightStatusTable
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/flights/airport/AirportMap
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /splitbookingflightreservation
Disallow: /splitbookinghotelreservation
Disallow: /rentals/
Disallow: /global
Disallow: /gmap
Disallow: /ugtm
Disallow: /gtm
Disallow: /mgtm
Disallow: /handlers/*
Disallow: /Handlers/*
Disallow: /QUkd4lO9/*
Disallow: /extra
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/search/seo
Disallow: /ugtm
Disallow: /search-widget
Disallow: /i/api/search/dynamic

User-agent: AdsBot-Google-Mobile
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /api/search/V8
Allow: /tweb/hotels/results-ajax
Allow: /tweb/hotel/history/
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /hotels/$
Allow: /hotels/*
Allow: /flights/$
Allow: /flights/*
Allow: /cars/$
Allow: /cars/*
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /sem/
Allow: /semi/
Allow: /in
Allow: /horizon/sem/
Allow: /*/landing/*.html
Allow: /tweb/hotels/
Allow: /tweb/flights/
Allow: /tweb/cars/
Allow: /charm/
Allow: /book
Allow: /s/tweb/session/refresh/presentation
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/flights/airport/AirportFlightStatusTable
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/flights/airport/AirportMap
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/flights/flightroutes/brands/momondo/DealsToCountryCities
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /splitbookingflightreservation
Disallow: /splitbookinghotelreservation
Disallow: /rentals/
Disallow: /global
Disallow: /gmap
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/search/seo
Disallow: /ugtm
Disallow: /search-widget
Disallow: /i/api/search/dynamic

User-agent: Google-HotelAdsVerifier
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /api/search/V8
Allow: /tweb/hotels/results-ajax
Allow: /tweb/hotel/history/
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /hotels/
Allow: /hotels/*
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /sem/
Allow: /semi/
Allow: /in
Allow: /horizon/sem/
Allow: /*/landing/*.html
Allow: /tweb/hotels/
Allow: /tweb/flights/
Allow: /tweb/cars/
Allow: /charm/
Allow: /book
Allow: /k/ident/
Allow: /s/ident/
Allow: /hotelreservation
Allow: /splitbookinghotelreservation
Allow: /mshotelreservation
Allow: /FDhotelreservation
Allow: /s/tweb/session/refresh/presentation
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /flights/
Disallow: /cars/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /carreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /splitbookingflightreservation
Disallow: /rentals/
Disallow: /gmap
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic

User-agent: Google-Travel-Flights
Allow: /book/flight
Allow: /flightreservation
Allow: /api/whisky/V5/flight/
Allow: /api/whisky/V1/userData
Allow: /api/pricePrediction/V1/flight
Allow: /api/moonshine/collect
Allow: /api/staticdata/whiskyStaticInfo/v1
Allow: /api/moonshine/V2/validatephone
Allow: /api/whisky/V1/flight/seatmaps
Allow: /api/whisky/V5/ack
Allow: /api/whisky/V5/error
Allow: /api/whisky/V1/abandon
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /flights/$
Allow: /hotels/$
Allow: /cars/$
Allow: /trains/$
Allow: /trips/users/
Allow: /cruises/$
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /charm/g/
Allow: /tweb/app/
Allow: /s/horizon/compareTo
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /flights/
Allow: /SNflightreservation
Allow: /msflightreservation
Allow: /FDflightreservation
Allow: /splitbookingflightreservation
Allow: /book
Allow: /in
Allow: /s/tweb/session/refresh/presentation
Disallow: /api/search/V8
Disallow: /tweb/hotels/results-ajax
Disallow: /tweb/hotel/history/
Disallow: /i/api/search/v1/hotels/poll
Disallow: /charm/horizon/cars/citycars/CityCarsAgencyMapViewLink
Disallow: /charm/horizon/cars/airportcars/AirportCarsResults
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /s/horizon/common/layout/StyleJamNavMenu
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/flights/flightdeals/frontdoor/FlightDealsLinks
Disallow: /charm/horizon/common/compareto/slide/SlideCompareToAction
Disallow: /charm/horizon/common/layout/MoreNavContentApiAction
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/flightroutes/AjaxGoodToKnow
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/flights/flightroutes/AjaxWhenToBookCharts
Disallow: /charm/horizon/flights/flightroutes/AjaxFlightRouteInfoTable
Disallow: /charm/horizon/flights/flightroutes/CountryCityRouteFAQAction
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/common/upgrade/UpgradeBrowser
Disallow: /charm/horizon/flights/airport/AirportFlightStatusTable
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /s/horizon/common/corporate/PlatformToBusiness
Disallow: /charm/horizon/cars/citycars/CityCarsAgencyMap
Disallow: /charm/horizon/flights/airport/AirportMap
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /vs/
Disallow: /%20/
Disallow: /maps/
Disallow: /tweb/
Disallow: /sem/
Disallow: /horizon/sem/
Disallow: /*/landing/*.html
Disallow: /semi/
Disallow: /hotels/
Disallow: /cars/
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /mscarreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDhotelreservation
Disallow: /splitbookinghotelreservation
Disallow: /rentals/
Disallow: /global
Disallow: /trains/
Disallow: /cruises/
Disallow: /car-static-data-requirements
Disallow: /restaurant-static-data-requirements
Disallow: /static-data-requirements
Disallow: /huddle/
Disallow: /guides/u/*
Disallow: /guides/admin*
Disallow: /guides/missing
Disallow: /guides/noaccess
Disallow: /s/horizon/common/personalization/guidebooks/
Disallow: /restaurants/
Disallow: /ugtm
Disallow: /curated/
Disallow: /nearby/
Disallow: /platform2business
Disallow: /playground
Disallow: /sandbox
Disallow: /benchmark
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic

User-agent: Mediapartners-Google
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /api/search/V8
Allow: /tweb/hotels/results-ajax
Allow: /tweb/hotel/history/
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /hotels/$
Allow: /hotels/*
Allow: /flights/$
Allow: /cars/$
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /sem/
Allow: /semi/
Allow: /in
Allow: /horizon/sem/
Allow: /*/landing/*.html
Allow: /tweb/hotels/
Allow: /tweb/flights/
Allow: /tweb/cars/
Allow: /charm/
Allow: /book
Allow: /s/tweb/session/refresh/presentation
Disallow: /hotels/
Disallow: /flights/
Disallow: /cars/
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/flights/airport/AirportFlightStatusTable
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/flights/airport/AirportMap
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /h/
Disallow: /s/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /labs
Disallow: /carreservation
Disallow: /hotelreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /mshotelreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /FDhotelreservation
Disallow: /splitbookingflightreservation
Disallow: /splitbookinghotelreservation
Disallow: /rentals/
Disallow: /gmap
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic

User-agent: AdIdxBot
Allow: /k/authajax
Allow: /h/mobileapis/
Allow: /f/smarty
Allow: /s/mobileutil
Allow: /api/search/V8
Allow: /tweb/hotels/results-ajax
Allow: /tweb/hotel/history/
Allow: /api/search/V8/hotel/
Allow: /i/api/search/v1/hotels/poll
Allow: /s/tweb/session/refresh
Allow: /h/xplanding
Allow: /hotels/
Allow: /hotels/sitemap
Allow: /cars/sitemap
Allow: /sem/
Allow: /semi/
Allow: /in
Allow: /horizon/sem/
Allow: /*/landing/*.html
Allow: /tweb/hotels/
Allow: /tweb/flights/
Allow: /tweb/cars/
Allow: /charm/
Allow: /book
Allow: /hotelreservation
Allow: /splitbookinghotelreservation
Allow: /mshotelreservation
Allow: /FDhotelreservation
Allow: /k/ident/
Allow: /s/ident/
Disallow: /charm/horizon/common/search/PreloadAction
Disallow: /s/horizon/common/layout/AjaxFooterLinks
Disallow: /charm/horizon/common/layout/AjaxFooterLinks
Disallow: /s/horizon/common/privacy/AjaxHeaderCookiesMessage
Disallow: /s/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/privacy/AjaxStyleJamHeaderCookiesMessage
Disallow: /charm/horizon/common/layout/NavMenuContent
Disallow: /charm/horizon/flights/cabinclassflightroutes/AjaxCabinClassFlightRoutesGoodToKnow
Disallow: /charm/horizon/restaurants/static_details/ajax/RestaurantDetailsReviewsList
Disallow: /charm/horizon/hotels/cityguides/CityGuidesBacklinkActivityUrls
Disallow: /charm/horizon/hotels/venue/ConventionCenterCarsResults
Disallow: /charm/horizon/flights/airport/AirportFlightStatusTable
Disallow: /charm/horizon/common/core/AjaxMany
Disallow: /charm/horizon/flights/flightroutes/LatestFlightDealsAjax
Disallow: /charm/horizon/flights/flightroutes/IpOriginAjax
Disallow: /charm/horizon/flights/airport/AirportMap
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /flights/
Disallow: /cars/
Disallow: /k/
Disallow: /r/
Disallow: /out
Disallow: /tracking
Disallow: /akamai-sureroute-test-object.html
Disallow: /mail/termsandconditions
Disallow: /clickthrough.jsp
Disallow: /empty.html
Disallow: /moira/
Disallow: /adclick
Disallow: /bookings
Disallow: /carreservation
Disallow: /flightreservation
Disallow: /mscarreservation
Disallow: /SNflightreservation
Disallow: /msflightreservation
Disallow: /FDcarreservation
Disallow: /FDflightreservation
Disallow: /splitbookingflightreservation
Disallow: /rentals/
Disallow: /gmap
Disallow: /charm/horizon/uiapi/
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/search/seo
Disallow: /i/api/search/dynamic

User-agent: BUbiNG
Disallow: /

User-agent: proximic
Disallow: /

User-agent: A6-Indexer/1.0
Disallow: /

User-agent: ADmantX Platform Semantic Analyzer
Disallow: /

User-agent: ContextAd Bot
Disallow: /

User-agent: berlin-fu-cow
Disallow: /

User-agent: ias-ir
Disallow: /

User-agent: ias-sg
Disallow: /

User-agent: *
Disallow: /charm/horizon/common/authentication/providers/AuthStateProviderAction
Disallow: /charm/horizon/react/component/PrivacyMenuStateProviderAction
Disallow: /charm/horizon/common/privacy/providers/CookiesDataProvider
Disallow: /charm/horizon/react/component/FooterBrandsStateProviderAction
Disallow: /charm/horizon/react/component/CompareToConfigStateProviderAction
Disallow: /search-widget
Disallow: /a/api/flightPricePrediction
Disallow: /tracker/

User-agent: AhrefsBot
Disallow: /i/api/seo/
Disallow: /i/api/hotels/image/v1/thumbnailsUrls
Disallow: /i/api/trips/
Disallow: /i/api/

Sitemap: https://www.kayak.com.sv/sitemap.xml
