User-agent: *
Disallow: /update/
Disallow: /install/
Disallow: /admin.php
Disallow: /admin/
Disallow: /config.php
Disallow: /license.html
Disallow: /readme.md
Sitemap: https://santillana.com.sv/sitemap

